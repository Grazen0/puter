`ifndef PUTER_CPU_IMM_EXTEND_VH
`define PUTER_CPU_IMM_EXTEND_VH

`define IMM_SRC_I 3'd0
`define IMM_SRC_S 3'd1
`define IMM_SRC_B 3'd2
`define IMM_SRC_U 3'd3
`define IMM_SRC_J 3'd4

`endif
