`ifndef PUTER_CPU_CSR_FILE_VH
`define PUTER_CPU_CSR_FILE_VH

`define CSR_MTVEC 12'h305
`define CSR_MEPC 12'h341
`define CSR_MCYCLE 12'hB00

`endif
