`ifndef PUTER_CPU_H
`define PUTER_CPU_H

`endif
